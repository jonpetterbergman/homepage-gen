Axis sv
