Axis
Axis min arbetsgivare
