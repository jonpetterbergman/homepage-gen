<navgen>
  <title>Ingen översättning hittades för denna sida</title>
  <content>
    <p>Ingen svensk översättning hittades för denna sida</p>
  </content>
</navgen>    
