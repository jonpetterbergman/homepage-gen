<navgen>
  <title>Axis</title>
  <content>
    <p>Axis min arbetsgivare</p>
  </content>
</navgen>    
