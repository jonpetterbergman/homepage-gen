<navgen>
  <title>Jobb</title>
  <content>
    <p>Blah Blah Jobb</p>
  </content>
</navgen>    
