Haskell
Haskell min hobby
