Jobb
Blah Blah Jobb
