<navgen>
  <title>Haskell</title>
  <content>
    <p>Haskell min hobby</p>
  </content>
</navgen>    
