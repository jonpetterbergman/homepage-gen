Hemsida
Petter Bergmans hemsida
