<navgen>
  <title>Hemsida</title>
  <content>
    <p>Petter Bergmans hemsida</p>
  </content>
</navgen>
